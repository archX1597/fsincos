class c_1397_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1397_2;
    c_1397_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz1z1x01x101x01zx1100z10z1xx01zxzzzzzxzxxxzzxxzxxzzzxxxxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
