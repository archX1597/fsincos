class c_1292_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1292_2;
    c_1292_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz110x1xx0xxzzzzzx1x100z0xz1zz0xxxzxxxxzzxzxzzxzzzxzzxzxzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
