class c_1092_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1092_2;
    c_1092_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzxx11011x011zx1x0xzxxz1x0x1xx0xxzxzzxxzxxxzxxxzxxzzzxxzzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
