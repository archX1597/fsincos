class c_1865_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1865_2;
    c_1865_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111z1xx0xz0xxxzx00zxz0111zzz1x1xxzxxxzxzxxzxzxxxzxzxxzxzzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
