class c_502_1;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_502_1;
    c_502_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1110z1z0xzx11110xxz1z0z0xx00z1xxxxxxzxxxxzxzxxzxzxxzxxxzzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
