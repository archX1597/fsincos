class c_1155_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1155_2;
    c_1155_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx0x0x00z1xzxxx1zxz1z111z01x00xzzxxxxzzzxxxxzzzxzzxzxxxxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
