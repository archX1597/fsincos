class c_1959_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1959_2;
    c_1959_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x001001zz1x1z00z100x01001xz0zzzzzzzxxxxzxzxxxzzzzzzxzxzzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
