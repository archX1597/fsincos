class c_1619_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1619_2;
    c_1619_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x01x0z0x1001x1zx0x110x100xxxz1zzzxxxzzxxxxzxzzxxxxxxxzxxzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
