class c_1708_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1708_2;
    c_1708_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111x0z1zz0zzx0xxz01001xz1x11z0z1zzzzxzxxzzzzxxzzxzzxzxzxxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
