class c_1989_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1989_2;
    c_1989_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z100x00zzz11z0xx010xx1x01xxx1011zxxzxxzxzzxxxxzzzzxxzzzzxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
