class c_1868_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1868_2;
    c_1868_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01101x0x0z01x011xz110xz1xx1zxzxxzxxzzxzxzzxzxxxzxzxxxzxzxxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
