class c_1434_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1434_2;
    c_1434_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxz110zx1x0xxz1x0xzzx0xzz000zx0xzzzzzzzzzzzxxxxxzxxxxzzzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
