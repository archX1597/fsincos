class c_1950_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1950_2;
    c_1950_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1z00001x10z1x1xxzzz11z110x1xzxzzxxxzzzzxzxxzzzxxxxzzzxzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
