class c_1587_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1587_2;
    c_1587_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110zxzzxxzzzz1x010z011zx1z00x1z1zxxzzxxxxxzzzzxxzxxxzxzxzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
