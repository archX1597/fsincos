class c_1732_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1732_2;
    c_1732_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx11x0x0x10z011101z0zx1001x1zz0zxzzzxxxzxzxxzxzxzxzxzzxzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
