class c_1588_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1588_2;
    c_1588_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10xz0z100zzxzzxzx1111zzx1z10111xxzxxxxxzzxxxxxxxxxzzzzxzzzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
