class c_1135_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1135_2;
    c_1135_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101xzxxxz01x10z1x1zzzzx1x0z1x0z0zzxxzxzxzxxzxzzxxxxxzxzzzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
