class c_312_1;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_312_1;
    c_312_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x00x1x1zxx10x011zx0z0zx1zz111x1xxxxzxxxxzzzzzxxxzxzzxxxzzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
