class c_1040_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1040_2;
    c_1040_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x011z1xz00zx000x0101zx10zz00xzxzzzxxxzzxxxzxxzxzzzxxxxzzxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
