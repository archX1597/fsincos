class c_1809_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1809_2;
    c_1809_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1x010101xxx10x1z0x0100x0zx11z0zzxxxzxzxxxzxxxxxxzzzzzzxzxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
