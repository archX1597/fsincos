class c_1966_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1966_2;
    c_1966_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1000zz00z10xzx0xx0x01xzzz0z0x0z1xxxxzxzzxxxxzxxxzxzzxxxzzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
