class c_1195_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1195_2;
    c_1195_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xxzz000zxzx1x0zzz01001xxzxz1zxzxzxzxxzzzxzzzzxxzxzxxzzxzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
