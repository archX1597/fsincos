class c_1663_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1663_2;
    c_1663_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1zx011x1zxxz0z100z0z0000zz00x0xzxxxxzzxxxxzxxxxxzzxzzzzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
