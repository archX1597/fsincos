class c_1272_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1272_2;
    c_1272_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0x0zx1x101z1100x000z0xzzzxx110zzxzxxxxxxxxzxxxzzxzzxxxxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
