class c_1496_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1496_2;
    c_1496_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxx01xzzz1z0z00x0z000xxz01zx01zzzxzxxzzzzzxxzzzzzxxzzzxzxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
