class c_1473_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1473_2;
    c_1473_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00111xz0zz1zzzz0z10zzx100x11x1zzzxzzzzxxzxxzxzxxxzzxzxxzzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
