class c_1540_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1540_2;
    c_1540_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100z110z0z11z11x01z0xxz1xxxxzxxzzxxxxxxzzzzzxxzxxzzxzxzxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
