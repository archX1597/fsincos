class c_1873_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1873_2;
    c_1873_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00010xzzx0z1zzx010zxxxx0xz00z0z1zzxzzxzzxzzxzxzzxzzxxzxzxzzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
