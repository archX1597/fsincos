class c_1896_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1896_2;
    c_1896_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzx00z001x11x01xx1z00xz101zzz01xzzzzxzzxzzxzzzzxxzzxzxzxxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
