class c_1974_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1974_2;
    c_1974_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1x0xzxx1x0zxz0000zx111xx000zxxxzxxxzxzzzzxxzxzxxzzxzzxxzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
