class c_1818_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1818_2;
    c_1818_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00xxzx1xz100x11xx0x10x0x0zxx0x0zxxxxzxxxxzxzxzzxxzxxxxzxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
