class c_1213_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1213_2;
    c_1213_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx101zxzzzx01zz001x1111zx1x01zxxzzzzxzzzzzxzzxzxzxzxzzzxxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
