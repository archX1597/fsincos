class c_1207_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1207_2;
    c_1207_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x011zzx10zx0x110zzxz01x0zx110x0xxzzzzzxxzxzzxxzxxzzzzzxzxxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
