class c_1594_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1594_2;
    c_1594_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111zz001xz0110z1011zx0zz0z001111zzzzxxxzxzxzxzxxxzzxxzxzzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
