class c_1767_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1767_2;
    c_1767_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z011xz1zxxzz01x1z10xxx000zx10x0xzzxzxxxxxxzzzxzzxzxxzzxzzzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
