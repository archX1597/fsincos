class c_1142_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1142_2;
    c_1142_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx10z01x11zx0xx01z111x0xzxzzx11xzxxzxxzxzzzxxxzxzzxxxzzxzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
