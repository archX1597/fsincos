class c_1574_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1574_2;
    c_1574_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzxzzzzz110x0z01zxz0zzx0zzzzz01zzxzzzxzxxzzzzxxxxzzzzxzzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
