class c_1278_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1278_2;
    c_1278_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x11zx000zx00x0111xz1z011zzx0xzxzxzxxxxxzzxzzzzxzxxzxxxxzxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
