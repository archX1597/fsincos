class c_1584_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1584_2;
    c_1584_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0x00zx1xz0zx0z110zx1x0zzx01zzzxzxxxzzzxzxxzzxzxxxzxzzzxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
