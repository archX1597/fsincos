class c_1837_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1837_2;
    c_1837_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzx0x1110z00x000x00zxxxx1z0z00xxzxzxxxzxzxxxxxzzzxzxxzzzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
