class c_1309_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1309_2;
    c_1309_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxz00z1x0x100110z00x0z1z1z1zz00xzxxxzxxzxxzxzxzxxxxxxzzxzzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
