class c_1652_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1652_2;
    c_1652_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xzz110111xz1xx010zx00xzzx0zxx0xzzzzzzxxzxzzxzzxxxxxxzzzxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
