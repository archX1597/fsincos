class c_1824_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1824_2;
    c_1824_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxzz0x1xx0x01zz0z01xz1zxzz1z00zzxzzxzxxzzzxzzzzzxzzxzxxzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
