class c_1237_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1237_2;
    c_1237_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz000x10zzxx1xxz10z1z01011x1zx1zzzzzxzxxzzxxxxzzxxzxxzxxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
