class c_1683_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1683_2;
    c_1683_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xz1xz11zx1x011xz01z1zz110x0x00zxxxzxzzxxzxxzzzzzzxxxxzxxxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
