class c_979_1;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_979_1;
    c_979_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z10x111zx10zx1z1zx00x1z0xx001x0xxzxxxzzxzxxzzxxxxzxzzxzxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
