class c_1263_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1263_2;
    c_1263_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0x0z01zx1zx1xz1x1x0zx00zz1x010zzxxxzxzzzxxzxxxxxxzzzzxxxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
