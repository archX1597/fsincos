class c_1382_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1382_2;
    c_1382_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10xxzxx1xzzx1101000111100x10z1xxzxxxzxxxxxzxxxxxxxzxzxxzxxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
