class c_1984_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1984_2;
    c_1984_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010x1zx111zz0101z001xx1x0xx01000zxxxzxxxxzxzzxxxxxxxzxzzxzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
