class c_1083_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1083_2;
    c_1083_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z11xx01z0xzz10xzzxzz00zx0xx0xzxxzxzxxzzxxzxxzxzzxzzzxxzxzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
