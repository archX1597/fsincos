class c_1122_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1122_2;
    c_1122_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xzx0x00zzzz0000zxx1zx01zx00x10zzxxxxzxzxzxxzxzzxzxxzxzxxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
