class c_1154_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1154_2;
    c_1154_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z111110zxzx01x0zz1z00x01xzz1zxzxzxxxzzzxxzxzzxzxzxzxzzzzxzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
