class c_1850_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1850_2;
    c_1850_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01011zz00x110x1z101x10z0x10zxxzzxzxzzzxxzxzxzxzzzzzxxzzzxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
