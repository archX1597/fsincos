class c_1688_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1688_2;
    c_1688_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zxxxz0001z1101xzx0111x111zz1zxzxzxzzxzzxxxxzzzzxxzzzxzzxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
