class c_1394_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1394_2;
    c_1394_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011z101xx00z0zz110x0x1xxz01zzzxzzzxxzxzzzzzzzzxxzxzzxzzxzxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
