class c_1291_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1291_2;
    c_1291_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1xzxx001x001zz00zz1z1zx111xx0zxzzzxzxxxzzxzzxxxxzzzzxzzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
