class c_1381_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1381_2;
    c_1381_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1x01zzx1zzz00x1x1001xx1x1001x1xzzxxxxzzxxxxxzzzxzxxzxzzxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
