class c_1998_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1998_2;
    c_1998_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1x10zxzxzz10z10z0x00xxx0zzz011xzxxxxxxxxxxzxxxzzzzzxxxxzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
