class c_1893_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1893_2;
    c_1893_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111010110xzzxz111zz00zx1xz10x0x1zzzxxxzxzzzxzxxxzzzzzxzxzzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
