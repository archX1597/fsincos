class c_1592_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1592_2;
    c_1592_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01x1zzz010x01zzxxz1zx111xx10x0xxxzxzxxxzxxzzzzzzxxxzxxzzzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
