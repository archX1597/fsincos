class c_1459_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1459_2;
    c_1459_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz11z0x01xx0xz00101xz0xx01111xzzzzzzzxzzzzzzzzxxzxxxxzxzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
