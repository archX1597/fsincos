class c_1672_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1672_2;
    c_1672_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0x0z11xzzx1x101z1x01x01z0zzz0xzxxxxxxzzxzzzxxxzzxxxzzxxxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
