class c_1164_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1164_2;
    c_1164_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x101zx0x1z0z00x1zz0x00z01zzzx1zzzxxxxzzzzzxxxxxzzxxxzxzzxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
