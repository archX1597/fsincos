class c_1464_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1464_2;
    c_1464_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zzz1zzzx1z11xxx0z00z01z1zz1x01zzxzzxzzzxzxzxxzzxxxxxxzzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
