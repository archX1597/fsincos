class c_1118_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1118_2;
    c_1118_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx0xx000010z1xx11zxxz1xxz0100zzxzxzxxxzzxzzzxzzzxxzxxxzzxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
