class c_1114_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1114_2;
    c_1114_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0xzx0zzxxzz1x0x0100z11zxz1zx1xxzzzxzzxxzxxxxzxxzxzzxzzxzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
