class c_1991_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1991_2;
    c_1991_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1x0xxz10xzxxxz11z110x1000x00z1zxxzxzxxzzzxzzzzxzxxzxzxxzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
