class c_1316_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1316_2;
    c_1316_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xxxx0z1z1z00zzxz10zzzx1z1zz1xxzxzzxxxzzxxzxzxxxzzxxxzxzzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
