class c_1902_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1902_2;
    c_1902_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zx10xzx11z0zxxz00xxz1zzzz00z01xzzxzzxzxxxzxzzxxxzxzzxzzzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
