class c_1999_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1999_2;
    c_1999_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx11z1xz0z001z1xxz00xz01z1x10zzxzzxzzxzzxxxxxxzxxxxzzzzzxzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
