class c_1117_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1117_2;
    c_1117_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx001010100z000xxxzzx010z1z00xzzzxzzxzxxzxzxzxxxxxxxxzzzxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
