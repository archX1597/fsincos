class c_1436_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1436_2;
    c_1436_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0xx0101x01zx1xx0x11x1001100zzxxzxzxxxzzxxzzzzxzzxxxzzzzxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
