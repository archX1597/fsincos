class c_1293_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1293_2;
    c_1293_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10x10z1z0xz100x0101z0xx11xz1000xzxxxxzzxzxzzxzxxzxzxzxzzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
