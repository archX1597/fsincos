class c_1611_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1611_2;
    c_1611_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10101zz0x0xxx11xx11zx0x00x1z0x1zxzxxzxzzxxzxxzzxxxxxzzzxxzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
