class c_1395_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1395_2;
    c_1395_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z0x01xx0z0zx0zx1x10x11xzxxxxx1xzzzzxxzzxzzzxxzzxzzxzzxxxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
