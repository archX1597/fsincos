class c_1607_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1607_2;
    c_1607_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx0z00z0111011zx00x0x1xxzz100zzzxxzxzxxzxxxxxxzzzxxzxzxzxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
