class c_1765_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1765_2;
    c_1765_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzx10zx00x0z0xx0x0x1xzzz01zxx00xzzzzzzxxxxzxxxxxxzzzzxxzxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
