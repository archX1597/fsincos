class c_1168_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1168_2;
    c_1168_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11zzx1z1x0z1100x0xz111z1xzxz1z0zxzxxxxxxzxxxxzzxxxzzzzxzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
