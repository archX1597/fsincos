class c_1658_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1658_2;
    c_1658_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz01z1xzz1x0z1x0z1z1zzxxz0z0xz0zzzxzxzzzxxzzzxzzzxzxxzxxxxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
