class c_1659_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1659_2;
    c_1659_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11001z10zxz01x11x11000z1xzz0110zzxxzzxxxzzxzxzxzzzxzxxxxxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
