class c_1371_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1371_2;
    c_1371_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10x00z0xz100100xxzzxx0zz1x1xzxz0xzzxxxzxxzzxxxxxzxxzxxxxxzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
