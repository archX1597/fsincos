class c_1129_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1129_2;
    c_1129_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zx110zxz10x0011x0zxx1xzz1z0x01xzzxzzzxzxxzzzzzzzxzzxxzxxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
