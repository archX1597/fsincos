class c_1079_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1079_2;
    c_1079_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx1zzx10x11x111xx0xz101z111zx01zzxxxzxzxxzzzxzxzzzzzzxxzxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
