class c_1687_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1687_2;
    c_1687_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx0z101xz0x10xzz10xz1zzz11z0zx0zzxxxxzxzxzzxzxzzzzxxxzzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
