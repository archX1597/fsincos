class c_1096_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1096_2;
    c_1096_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0110x10zz1xzzz1zz00z1zxzz11xxzzzzxzxxzzxzzxxzzzzxxxzzxzzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
