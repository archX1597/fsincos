class c_1286_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1286_2;
    c_1286_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z0z1x10x1x0x1xxx01x0x11z00010zzzzxzzxxxxzxxxzzzxzzzzxxxxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
