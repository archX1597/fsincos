class c_1962_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1962_2;
    c_1962_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z01z00001xz1010xz0zxzz0xzz110xxzzzxzzzxzxzxxzzzxzzzxxzzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
