class c_1105_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1105_2;
    c_1105_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11zx1x00xx0z010xxxz00x11zz0zxxzzzxxxxxzxzxzzzxxzxxzxxxzzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
