class c_1072_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1072_2;
    c_1072_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00000x10100z1z1xxz0z0zxxz00x0z1zzzzxzxxzzzxzzzzzzzxxzxzzzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
