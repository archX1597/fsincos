class c_1485_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1485_2;
    c_1485_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z01xz10zx0z1x1011z11zz101xxzx1zxzzxxzxzxzxxxxzzzzzzxxxxzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
