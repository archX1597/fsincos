class c_1859_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1859_2;
    c_1859_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx101x1z0xxzx00x1z00110zx0x1xz0xxzzxzzzxxzzxxxzzxxzxxzxzzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
