class c_1564_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1564_2;
    c_1564_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx11zxxzz0xxx1x1zx10xzxz1xx1xz0zxzzxzzxzzzzzzxxxzzzxzxzxzzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
