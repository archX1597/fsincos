class c_1167_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1167_2;
    c_1167_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0x1zx0zxx0001z01xxzzxxz1xx11x0zxzzzxxzxxxzzzzzxzzxzzxxxxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
