class c_1311_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1311_2;
    c_1311_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1z1z0z1x00z00zz10x10x01001zz0zxxxzxzzzzzzzxzzxzxzzzzxxzxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
