class c_1774_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1774_2;
    c_1774_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z11xxz11x01zzx0000xzx1z11x011xzzxxzzzxxxxxzzxzxxxzzzzxzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
