class c_1783_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1783_2;
    c_1783_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0z111x110zx10x0x01010zx1xz0xzzzxzzxzzxxxxzzxxzxzxzxxxzxxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
