class c_1479_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1479_2;
    c_1479_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzz01x1x011x01zzxxxx1z1xzxxxz11xxxxxxzzzzxzzzzzxzxxzxzzxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
