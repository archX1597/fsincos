class c_1835_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1835_2;
    c_1835_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1101z1xx00zz0xxzz10xx010zxxz0z0zzzxzzxzxzzxzzxxzxxxxzzzzxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
