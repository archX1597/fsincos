class c_1268_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1268_2;
    c_1268_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0z1xzx001011001z0zz0zxxz11zx1zzzxzxxzzxxxzxxxxzxxxzxzzxzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
