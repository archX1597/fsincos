class c_1971_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1971_2;
    c_1971_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00x11zxx00xz0zz0xzxz01xz10xz0x1zxxzzxxxxxxxxxzzxzxxxxxxzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
