class c_1415_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1415_2;
    c_1415_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1100z01101xx10x00zz0zx0x0x1z0z0zxzzxzxzzxxzzzzzzxzxxzxzxxxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
