class c_1190_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1190_2;
    c_1190_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1x010xzzzx110xzx10z11xxz01x000zxzzxxzzzzzzxxxxxzxxzxzzxxxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
