class c_1449_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1449_2;
    c_1449_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzz10z10001zz0z11z00x0xx110x10xxxzzxxzzxxxxzzzzzxxzzxzzxzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
