class c_1789_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1789_2;
    c_1789_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z1z11zx0zz0x11x1zzzz1xz010z1zxzxxxzxxxzxzzzxzxxxzzxzxxxzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
