class c_1296_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1296_2;
    c_1296_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxx0xz10z00xxxxzx1001zx1x1z00xx0zzxzzxzxxzxzzxxxzzxzxxzzxzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
