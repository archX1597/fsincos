class c_1787_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1787_2;
    c_1787_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzz0z0z011xz0x0xzxxxx0zz000z10zzzxxxzxxxxzzxzzxzxxzxxxzxzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
