class c_1562_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1562_2;
    c_1562_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000xzx0011010z101110x01z11x1x1x0zzzxxzzzxxxzzxzxxzxzzzzzzzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
