class c_1954_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1954_2;
    c_1954_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xz11z10zx100x10x110x010x101z11xzxzxxxzxzzzzzzxzzxzzzzzxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
