class c_1466_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1466_2;
    c_1466_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x110zx1xx00zz1x1x0z1x1z0x11x00zzxzxxzzxxxzzxzzxxxxzzxzzxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
