class c_1196_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1196_2;
    c_1196_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xz011x0zxzxz0zxzx011z00x1zz0xzxxxzxxxxxzzxxxzzxzzzzxzxzxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
