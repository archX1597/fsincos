class c_1689_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1689_2;
    c_1689_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxzx10z11z0zzxx0x1x0xx010x1zx00zxzxzzxxxxzzxzxzzxxzzzxzzxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
