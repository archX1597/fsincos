class c_2001_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_2001_2;
    c_2001_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1111xzzx010001011z1zxz0xz001x1zxxxzxzzxzxzxxzxxzzzzzxxzzxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
