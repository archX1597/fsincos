class c_1341_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1341_2;
    c_1341_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1000x00110110xx0zzx01xx1x111z1xxxzxxxzxxxzxzxzzzzxxxzzxzxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
