class c_1613_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1613_2;
    c_1613_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01010101001x1111zxxzz0x00zzx0x1xxxzxzzxxzxxxxzxxxzzzzzxzxzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
