class c_1575_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1575_2;
    c_1575_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z10zz000xz101zzzz1z1x1zxx01z00xzxxzxzxzzzxxxzzxzzzxzxxzxxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
