class c_1534_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1534_2;
    c_1534_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zz010zxz0xzz10xxz01x1xxzz0010zzxxzzzzzxzzxzxzzxxxzxzzzzxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
