class c_1351_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1351_2;
    c_1351_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z1zzz1x0010x11x0x0z1xxz01xz0xxzzxzzxzxxzxxxxxzxxxxxzzxxzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
