class c_1208_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1208_2;
    c_1208_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1111z00xxzx0zx101z001zzzxzz111zxzzxxxzxxxzxzxxzzxzzxzxxxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
