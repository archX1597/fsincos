class c_1798_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1798_2;
    c_1798_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111zx1zxzx0zxxxzz0010zz0z11xzzzzzzzzxxxzzxzxxxxxzzzzxzzzzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
