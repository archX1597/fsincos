class c_1601_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1601_2;
    c_1601_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110x1000xxxxxzxxx0011x1zz110z0z1xxzzzxxxzxzzxxzxxxxzxzzxzzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
