class c_1784_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1784_2;
    c_1784_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0101x0z00xxz011x01z0x1x1x011z0x1xzxxxzxxzxzxzxxxzxzxzxzxzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
