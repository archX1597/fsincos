class c_1509_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1509_2;
    c_1509_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxzz1zx11x011x0x111100x01xz1zx1xxzxzxzxxzzxxzxzxzxxzxxxzxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
