class c_1786_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1786_2;
    c_1786_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxz1xxz10xzxx0z0zx01x11z0zz1zxzzzxxzzxxxzzxxzzxxzxxxxxxzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
