class c_819_1;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_819_1;
    c_819_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx000z110zzzz1z110x1zz0x10x11zxxzxxxxzzzxxxxxxzzxxzxzzzzzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
