class c_1323_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1323_2;
    c_1323_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z0xxxxzz0z110111zz10z1z1101z01xzzxzxxzxxxzxzzzxxzzzzxxzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
