class c_1532_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1532_2;
    c_1532_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxx1xzzxx011xx01x0z01x1100xxz00zxzzzxzxzxzzzxxzzzxzzxxxzzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
