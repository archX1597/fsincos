class c_1306_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1306_2;
    c_1306_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xx0xz01z0z1xz000z1x0000xx0101zzzxxzxxxzxzxzxzzxzxxxxxxzzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
