class c_1727_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1727_2;
    c_1727_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z0xz01zxz0xzzzz1x0x1z1z11x101xxzxxzxzxxxxxxzxxxzxxxzxxzxxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
