class c_1720_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1720_2;
    c_1720_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010zzx0zzxz1zzz1xxzz1z11101xzzxzxzzxzzzzzxzxzzzzxzzxzxxxxxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
