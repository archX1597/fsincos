class c_1770_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1770_2;
    c_1770_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1z0zx00zzz01x000zzzz01111x1xzxzzxxxzxzxzxzzzzzxxxxxxzxxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
