class c_1369_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1369_2;
    c_1369_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz101z01x1zzxzzxzzz1z1xxxzx01xxxxxxzxzxxxzzzxxxxzxzzzxzzzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
