class c_1474_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1474_2;
    c_1474_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx00zxz1110zxz00101z11x11011zz1zzxxzxzzxzzxxzxxxzxxxzzxzxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
