class c_1851_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1851_2;
    c_1851_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z0xxz1zz1111000z0zxz0xxxx0010zzzxzxxxxxzxxzxxxxzxzxxzzzxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
