class c_1953_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1953_2;
    c_1953_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz01xz0x1x0x1x10x1z1z010x101zz1zxzxzxxzxzxxzxxzxxxxxzzzzzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
