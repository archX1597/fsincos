class c_1322_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1322_2;
    c_1322_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101zxx0xzz0zx0zzzxxxx110z1z1z0z0zxzzxzzzxzzxzzzzxxzzxzxzzzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
