class c_1653_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1653_2;
    c_1653_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00xxz11011zz0zz0xz1z1x1xx01zzxxxzxxzzxxxxxxxxzzzzzzxxzzxzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
