class c_1821_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1821_2;
    c_1821_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx0xx01x01000xx0zzx11x1zxx1z10zxzxxzzxzzzzzxzzxxxzzzxxxzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
