class c_1244_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1244_2;
    c_1244_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx1xxzzxxx0x1xz00zz11xzxx0101zxxxzzzxxxxxxxxxzzxzxzxxxxxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
