class c_1747_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1747_2;
    c_1747_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z111zx00zz11111x110111x0011z101xxxxzxzxzzxzzzxzxxzzzzxxzxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
