class c_1099_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1099_2;
    c_1099_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx00zzz0z1xx11x0x0x10x1x0xx11zxxxzzzzzzxzxxxxzzxxxzxxzxzxzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
