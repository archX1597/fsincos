class c_1606_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1606_2;
    c_1606_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z01z11101x101x11xz0x0zz0001x010zxxzxxzxzzxzxxxzzxxxzxzzzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
