class c_1163_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1163_2;
    c_1163_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzx1xzx10xzzzx0z1x10x01101zxx00zxxzzzzzzzzzzzzxzxzxxxxzxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
