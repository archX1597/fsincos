class c_1507_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1507_2;
    c_1507_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xx00xxx101x11z0xzz11x1z1zz111zzzxzzxzxzzxxzxzzxxzzzxxxzxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
