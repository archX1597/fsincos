class c_1945_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1945_2;
    c_1945_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx1z1xz101xz011z1x0zz11xz0zzz11zxxzxxxxxxxxzxxxxzzxzxzzzxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
