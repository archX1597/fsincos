class c_855_2;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_855_2;
    c_855_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z011z00x101x0zzxx01zzzxx1z1x01xzxzxzxzxxxzxxxzzxzxzxxzxxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
