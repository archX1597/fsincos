class c_1576_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1576_2;
    c_1576_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1zx0x01z0z1x1110x01z00xxx0x111xxzzxxxxzxzzxzzxzxxxzzzzxzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
