class c_1826_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1826_2;
    c_1826_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zzx1xx0x0z0xzzzz1x0xzzzx1xx0xxzzzzzzzxxzxxxzxxxzxxxzzzxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
