class c_1811_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1811_2;
    c_1811_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101zxxzzx10xxx10zx0zzxzxz0x1x1z1zzxxxzzzzxzzxxxzxxxxzxxxxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
