class c_1833_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1833_2;
    c_1833_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011x01110z110xxzxzzx0xz1000z0x1xxxxxxxzxzxxzzzxxzzzzxxxzxxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
