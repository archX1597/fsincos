class c_1234_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1234_2;
    c_1234_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z11x0z00zx0x0zxz0zxzz01xx0zzz1xzzxxzxxzxzzxzzxxxxxxxzzzxxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
