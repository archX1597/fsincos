class c_1313_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1313_2;
    c_1313_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzzz1zzz00x00zxz000xx1zzxz1zx10zxzxxzxxxxxxxxxzxzzzxzzzxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
