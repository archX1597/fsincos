class c_1214_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1214_2;
    c_1214_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x001xx1x1zz1101zx0x011zx01110x1xzxxzzxxzxzxzxxxzzxxxzxxzxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
