class c_1011_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1011_2;
    c_1011_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx11zx00z0x1xxzxz110x001z00zz111zxzzxxxxxzxzzxzzxzxxzzzxzxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
