class c_1808_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1808_2;
    c_1808_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz00x0xx00zzzz1zxzx0zxxzzz00xz0zxxzxzxzxxxzzxzxxzzxzzxzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
