class c_1503_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1503_2;
    c_1503_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1111x1x1000x11zz1xx010zz11x0z0x1zzzzxzzxxzzzxzzxxzzxxxzxxzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
