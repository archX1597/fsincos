class c_1201_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1201_2;
    c_1201_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxzzzxxzz1xz1xx001zz1xxzxxzx11xxxzzxzxxzxxxxxzzzzzxzzzxzxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
