class c_1982_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1982_2;
    c_1982_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz0xx101xxx00z0x10xxx1z011x00xzzzzzzzzxxzxzzzzzxxzxxxzxzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
