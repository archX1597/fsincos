class c_1726_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1726_2;
    c_1726_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzx0010z1xx0010110xzzx1xxz0x00zzxzxzzxxxxxzxzxzzxzxxzxxzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
