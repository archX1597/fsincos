class c_1895_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1895_2;
    c_1895_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100x0xz0x1xxzxx1xzzzzx0101x10111xxzzxzxxzxxzzzxxzxxzzxxzzzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
