class c_1052_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1052_2;
    c_1052_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1zz101z1z101z1z0x1zzz1zzzxz000zzxxxxxzxzzzxxzxxxxxzzzzxzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
