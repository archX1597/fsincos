class c_1064_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1064_2;
    c_1064_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx000010xzx1xz11x0z100z1x1z0xx0zxxxxxzxzxzxzzzxxxxzxzzxzzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
