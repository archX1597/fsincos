class c_1905_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1905_2;
    c_1905_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0zxx1xzx1zzzx11000zx00101x1xxxxzzxzxxzzzxxxzxxxxxzxzzzxzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
