class c_1723_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1723_2;
    c_1723_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zzxzzxxz1zz10x011z1zz0x00x1z11xxzzzxxzxxzxxzzxzzzzxxxxxxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
