class c_1433_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1433_2;
    c_1433_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00xx00xxz01zxx0z0xz00100xzzz0z1xzxxxzxzzxxxxzxzxxzxzxzxzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
