class c_1807_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1807_2;
    c_1807_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0101x0z0x0zz1z11zzx10x1z1xx010zxxxxzzzzxxzxzxxzxxxzxxzxzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
