class c_1968_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1968_2;
    c_1968_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1100xxz1xx11z1xxz1zxxzx01xzz0x0zzzxzzzzxzxzxxxxxxzzxzxzxxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
