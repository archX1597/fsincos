class c_1486_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1486_2;
    c_1486_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z1xzx11x1z0z010xxx0z101z0x1x10xxzzxzzzzxxxxzzxzxxxxzzxzzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
