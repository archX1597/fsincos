class c_1150_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1150_2;
    c_1150_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0011zz11000z000x00z01xx001101110zxxxxxzzzzzxzzzzzzzzzzxxzzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
