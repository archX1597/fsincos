class c_1517_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1517_2;
    c_1517_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxz0xzx11x010x10z0z111z0010x11xxzzxzxxzzzzxxxxxzzxzzxzzxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
