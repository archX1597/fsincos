class c_1677_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1677_2;
    c_1677_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zx0x1z010zxx000x0100z10z10z0zxzzzxzxxzzzzzxzxxxxzzzxzzxxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
