class c_1465_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1465_2;
    c_1465_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xxz0x10x1xxxzxx010z11xzzxxz0zx0xxxzzzzzzzxzzzzxxxxzzzxzzzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
