class c_1034_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1034_2;
    c_1034_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x00z01xz0z1zx1x001x01z0zzzzzx0zxzzzzxzxzzxxzxxxxxzxxxxzzzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
