class c_1108_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1108_2;
    c_1108_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010xxxx000xzxz11zx1x1z10xxz1x1x0zzzxzxzxxzzxxxxzxxzzzxxzxzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
