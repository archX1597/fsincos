class c_1518_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1518_2;
    c_1518_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11111xxzxx010zz0z011zzx1zxz1010xxzzzzzxxxxxzxzzzxxxzzzzzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
