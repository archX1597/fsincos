class c_1836_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1836_2;
    c_1836_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zz10010zxx01zx1z0z1z1z01xzzzz0zxzzxzzzxxxxzzzxzxzxxxxxxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
