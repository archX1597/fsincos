class c_1570_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1570_2;
    c_1570_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx0z0xzx0xz000zxx0xxx01zx000zx0xzzzzzzzzzzzxxzzzxxzxzxzxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
