class c_1691_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1691_2;
    c_1691_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx110z1xz1x0xx0xzzzxx0z1zx00zx1xxxxxzxzxzzxxzzzxzxxzzzzzzzzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
