class c_1558_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1558_2;
    c_1558_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xx0zzzxxx0z0z11x00x011xx1z101zzxxzzzzzxzzxxzxzxxzxzzxxxxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
