class c_1759_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1759_2;
    c_1759_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzx0xxxz10zx1xx000z1z01zzz1x01zzzxzxzxxxzzzxxxxxzxxxxxzzxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
