class c_802_1;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_802_1;
    c_802_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1110x10z0z0zzzzx0x0z1x1zx0zz1x1xxzxzxxzzxzxzxzxxzxxxzzzxzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
