class c_1429_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1429_2;
    c_1429_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz0zzx0xz111xxx11zxxzx110z10zx0zzzzxxxxzxxzzxxzxxzxzzxxzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
