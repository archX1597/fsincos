class c_1442_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1442_2;
    c_1442_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100zxx010x11x1xz100zz0z11x1x0x1zxxxzzzzzzxzzzxzxxzxxzxxxzxxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
