class c_187_2;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_187_2;
    c_187_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z110z00x0z01xxxx1z1zxz0x010zx1x1xzxzxzxxxxzxzxxzzzzzzxzzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
