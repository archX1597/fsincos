class c_1377_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1377_2;
    c_1377_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x001z00x1z00x110zxxzx10zz0zx1010zxxzxxzxxxzxzzxzzxzzxzxxxzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
