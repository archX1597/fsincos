class c_1560_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1560_2;
    c_1560_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxzz1010z01xx1zz0z0zx001xx00xx0xxzzzzzxzzxxzxzxzzzzxxxxxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
