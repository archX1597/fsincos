class c_1380_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1380_2;
    c_1380_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zxz0zz10zx01zz0x11x0zxz1zz1x00zxzxxxzzzxxxzxxxzxxxzxzxxxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
