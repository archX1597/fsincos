class c_1284_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1284_2;
    c_1284_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzz1x1x0z0100x10zzx1100z00z0xz0xzzzxxxxzxzxxzxxzzxxxxxxxxxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
