class c_1963_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1963_2;
    c_1963_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxx011zxx0x01x01x1zxxz1z000zz11zzxxxzxzxzzxzxzzzzxzxzxxxxxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
