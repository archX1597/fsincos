class c_1492_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1492_2;
    c_1492_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx0x0x0zx1zxzzz00x0001zz000z01zxxzxxxzxxxzxxxxzzzzzxzxzzzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
