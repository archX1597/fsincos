class c_1917_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1917_2;
    c_1917_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzz00x11x01101zzx0x1zz01zz110xxzzxzzzxxzxxzzxxxxxxzzzzxzzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
