class c_1502_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1502_2;
    c_1502_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01101x110x0xzzx1zzxxz0xx10x0001zzzxzxxzxzxxzzxzxzzxzzxxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
