class c_1515_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1515_2;
    c_1515_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1zzz1zx1101101z1x101x10x1x1xzxxzzzzzzxzzzzzzxzzzzxxxxzzxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
