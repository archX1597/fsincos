class c_1396_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1396_2;
    c_1396_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z101xxzz10x1101xz0zx01zx01z01x0zzxzxxzzxzxxxxxxzzzzzxxzxxzzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
