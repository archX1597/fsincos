class c_725_1;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_725_1;
    c_725_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1zx0x111z0z11z0zx01x000zxz11x1xzxzzzzxxzzzzzzzzzzxzzxxzzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
