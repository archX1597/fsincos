class c_1915_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1915_2;
    c_1915_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxzzzx11z0xxx010zxx11zzx0zz01xzxxxxzzzzxxzzxzxxxzxzxxzxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
