class c_395_2;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_395_2;
    c_395_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz11xxx1001x1111010x0zz0zx0xz001xzxxzxzzzxxxzxxzxzxxzzzxzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
