class c_1269_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1269_2;
    c_1269_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz0z00zxxxxx1xz0001xxz011001zz1zxxzxxxxzxxzxxxzzxzzxzzzzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
