class c_1847_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1847_2;
    c_1847_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzz0xxxxz1z10x100z0110100xz0xz0xxxzzzxzxzzzzxzzxzxzxxzzxzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
