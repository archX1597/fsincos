class c_1899_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1899_2;
    c_1899_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101z00110xx1x11101x0011zxx1z0x1zzxxxxzxzzzzxxxzxzxzzzxzxxzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
