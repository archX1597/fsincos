class c_1678_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1678_2;
    c_1678_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01z111zxz00zxxzz0xz0xxzxxx01x1xzzzzzzzzxzzxzzzzxxzzzzxxxxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
