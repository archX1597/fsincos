class c_1349_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1349_2;
    c_1349_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1xx0z1z11x0x11000xxz10z100x010xxzzxxxzxzzxzxzzxxxzzzzxzzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
