class c_1470_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1470_2;
    c_1470_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0x0001xzxx10x1zxz1x1z0010x01x1xxzxxxzxxzxxxxxxxzxzxzzxzzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
