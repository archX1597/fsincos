class c_1709_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1709_2;
    c_1709_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz0001zx1x00101zzz0zxx00001z01zxzxzxzxxxzxxzzzzxzxzzzzxzxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
