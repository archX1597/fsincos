class c_1252_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1252_2;
    c_1252_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxxx1xxz1xzxz1x100z001zx0xzx01zxxzzzzzzzzzxzxzxxxxzzxzzzxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
