class c_1339_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1339_2;
    c_1339_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzx0xx0z0zzz0x10xxzx11xx11z00zx0zxzzzxxzzxxxzzxxxxzxzxxxxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
