class c_1236_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1236_2;
    c_1236_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101zz1z0zz10x1zxzxzxxx011001x0z1xxzzxzzxzzxxxxxxxxxzxzzzzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
