class c_1140_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1140_2;
    c_1140_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010zzz0z101010x11101z10x11001101xxxxxzzzzxxzzzxzzzxxzxzxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
