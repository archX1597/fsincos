class c_1280_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1280_2;
    c_1280_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzzz00xz0111011x001xzx0z100xx01xxxxzzzxzzxxxzxxxzzxxxxxxzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
