class c_1980_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1980_2;
    c_1980_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzx11z1zx0xzz0zzxxx00z111x0x10zzxxzzzxxzzzxzzzxxzzxxxzxxxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
