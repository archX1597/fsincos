class c_1764_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1764_2;
    c_1764_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz1zzxxxx01zz0x000xz1z1xzxxx01zzxxzxxxxzxzzxxzxxxzzzzxzxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
