class c_1729_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1729_2;
    c_1729_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10011zzxx00x00011x0zz0z100z1101xxzxzxzxxxzxxzxzzzxzxzxzxzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
