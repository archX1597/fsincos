class c_1886_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1886_2;
    c_1886_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz10x1x00zxzxzz1110zx100z0zzz010zxxxzzzzxxzxxxxxxzxzxzxzxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
