class c_1211_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1211_2;
    c_1211_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0000xxxxx10xz0z1zzx0xx00xz0zzzzxzzxzzxxxzxxxxxxxxxzxxzxzxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
