class c_1825_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1825_2;
    c_1825_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz010x1z0zzx11xx001zxxzxx1xx11x0xxzxzzzzzzzzxzxzxzzzxzzxzzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
