class c_1020_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1020_2;
    c_1020_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz00xz0xz01x01zxx101xzzz1z000zzxzxzzxxzxzzxxxzxzxzxxxzzzzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
