class c_1861_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1861_2;
    c_1861_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z01x1z11x01xz011z10z1z1zzzx0zxxxxxzzxxxzzzxxzzxzzxzxzzzzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
