class c_1495_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1495_2;
    c_1495_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxx10zxx01x0zx01zx0001xzxz1z10xzzzxzxxxxzxxzzzzxzzxxxxxxzxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
