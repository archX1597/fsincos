class c_1445_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1445_2;
    c_1445_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10100z0000z1xz111zxx11x1101z1x1xxxzzxzzzxzxxxzzzzxxzxzxzzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
