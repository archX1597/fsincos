class c_1317_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1317_2;
    c_1317_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z01zx0z1xz11z1110z101xxx11xzx1xxzzxxzxzzzzzxxzxxzzxxxzxzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
