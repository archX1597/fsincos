class c_1546_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1546_2;
    c_1546_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzxxzz0xz000zx1zxxz00x1zxz1xx10xxxzxzzxzzzzzxzxzzxzzzzzxxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
