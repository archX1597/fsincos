class c_1049_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1049_2;
    c_1049_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10z010z1zxz0x001z0z1000x0011x1xzzxxxzxxzxzxzxxzzxxzxxzzzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
