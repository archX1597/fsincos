class c_166_2;
    rand bit[7:0] f41_exp8; // rand_mode = ON 

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (f41_exp8 == 8'hfc);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../UVM_ENV/f41_sequence.sv:14)
    {
       (f41_exp8 <= 8'h80);
    }
endclass

program p_166_2;
    c_166_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10xzx0xxzz0zz000xxxzx0xxz0xx1x01xxxzxzzzxzzxzzxxzzzzzxxzxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
