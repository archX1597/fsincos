class c_1892_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1892_2;
    c_1892_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x0000111z01x0x0zx000101z0z101xxxzzzxxzzzzxzzzxxxzxzxzxxzzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
