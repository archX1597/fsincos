class c_1782_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1782_2;
    c_1782_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0z001zz110zxx0111zzz00x1x011z1xxxxzxzxxzzzxzzzzzzzxxzxzzxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
