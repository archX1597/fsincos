class c_1578_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1578_2;
    c_1578_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz00z10xz01zxz10z011110zx01z01zxxxxzzzxzxxxxxxzzxzxzzxxxxxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
