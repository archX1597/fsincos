class c_1062_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1062_2;
    c_1062_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz011zz00x00zzz0zz0001zxzzx1xx1zxxzzxzzzzzzzzzxzxxxxzxzxxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
