class c_1361_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1361_2;
    c_1361_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x010x10z0101z10x01z1zzx0zxz10z0zxzzzzxzzzxzzxzzzzzzxzxxxxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
