class c_1920_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1920_2;
    c_1920_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzzxzx0x010x0xzz00xx00x1101x01xxxzxzxxxzzxzzxxzxzxxxxxzxxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
