class c_1359_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1359_2;
    c_1359_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zzz11x0x0zzz1000z1011z0x00x1zxzxxxzzxzzzzxxzzxzxzxzxzxxxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
