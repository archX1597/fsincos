class c_1404_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1404_2;
    c_1404_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxzz10000x1zz1z00z01x11x0z110zzzxzzzxxxzxxxzxxzzxxxzzxzzxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
