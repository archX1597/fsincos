class c_1329_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1329_2;
    c_1329_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzzxz0x0x0x1xz1z0zz0xxxzxz110xxzzzxzxzzzzxxxxxxxzxxxxzxxzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
