class c_1408_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1408_2;
    c_1408_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z1z1z01x010z00zx1zzzzx1xxxz1xxxxzzxxzxzxzxxxzzxzzzxxxzxzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
