class c_1889_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1889_2;
    c_1889_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz01x1zz00x00x1x1xxz010x0x00zz0xzzzxxxzzxzzzxzzzxxzzxzzxzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
