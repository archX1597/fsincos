class c_1703_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1703_2;
    c_1703_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00zzxzx10x10xx00000xz001z1x1111zzzxxxzxzzzxxzxzzxzzxxxzxzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
