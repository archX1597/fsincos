class c_1290_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1290_2;
    c_1290_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z11xzx1zz01zx101z0xzz0x0zz0z01xxzxzzxxxxxzzxzxxzxzxzzzxzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
