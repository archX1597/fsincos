class c_1874_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1874_2;
    c_1874_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx11z01110x0xxz110xx10011xxxz001zzxxzzzzzxzzxxxzxzxxzxzzzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
