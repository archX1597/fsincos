class c_1623_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1623_2;
    c_1623_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101x10100z1x1xx00zxz0010zzxzxxxzzxzxzzxzzxzzxzxzxzxzxxzxxzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
