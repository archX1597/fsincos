class c_1545_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1545_2;
    c_1545_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx0z0101x10x10111z01z011z10x11x1xxzzzzxzxxzxzzxxxzzzxzxxxxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
