class c_1247_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1247_2;
    c_1247_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00z0x0zxz010100x0zz0x0xzz1zx1z1xxxzzzzxzzzxxzzxzzxxxxzzxxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
