class c_1804_2;
    bit[31:0] frac32 = 32'h0;

    constraint cons_this    // (constraint_mode = ON) (../UVM_ENV/f_transaction.sv:29)
    {
       (frac32 > 32'h80000000);
    }
endclass

program p_1804_2;
    c_1804_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0z1zzz0x1zz100zxx1x101zzz1xz1xxxxxzxxzxxxxxzxzxzxxxxxxxxxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
